library verilog;
use verilog.vl_types.all;
entity vector_tb is
end vector_tb;
